architecture pmRX_a of pmRX_e is

begin


end pmRX_a;
